module ysyx_22050612_EXU(
input imm,
input opcode,

input Mr_val,
output Mr_addr

);



ysyx_22050612_RegisterFile #(ADDR_WIDTH = 5, DATA_WIDTH = 64)(

);








endmodule
