module ysyx_22050612_TRANSPOSED_MATRIX(
	input [131:0]p00,p01,p02,p03,p04,p05,p06,p07,p08,p09,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,
	output [32:0]o00,o01,o02,o03,o04,o05,o06,o07,o08,o09,
	             o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
                     o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,
                     o30,o31,o32,o33,o34,o35,o36,o37,o38,o39,
                     o40,o41,o42,o43,o44,o45,o46,o47,o48,o49,
                     o50,o51,o52,o53,o54,o55,o56,o57,o58,o59,
                     o60,o61,o62,o63,o64,o65,o66,o67,o68,o69,
                     o70,o71,o72,o73,o74,o75,o76,o77,o78,o79,
                     o80,o81,o82,o83,o84,o85,o86,o87,o88,o89,
                     o90,o91,o92,o93,o94,o95,o96,o97,o98,o99,
                     o100,o101,o102,o103,o104,o105,o106,o107,o108,o109,
                     o110,o111,o112,o113,o114,o115,o116,o117,o118,o119,
                     o120,o121,o122,o123,o124,o125,o126,o127,o128,o129,
                     o130,o131
	     )

assign o00 = {p00,p01,p02,p03,p04,p05,p06,p07,p08,p09,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,

generate
	for



endmodule
