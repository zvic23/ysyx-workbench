//import "DPI-C" function void ebreak ();
import "DPI-C" function void set_gpr_ptr(input logic [63:0] a []);

`define ysyx_22050612_rgsize 64

module ysyx_22050612_npc(
input clk,
input rst,

//output [31:0]inst,
output [63:0]pc,

output [63:0]wb_pc

);

wire [31:0]inst;
wire [63:0]dnpc;
wire pc_update;

wire [63:0]imm_I;
wire [63:0]imm_U;
wire [63:0]imm_J;
wire [63:0]imm_B;
wire [63:0]imm_S;
wire [ 5:0]shamt;
wire [ 4:0]rd;
wire [ 4:0]rs1;
wire [ 4:0]rs2;


wire exu_block;


assign wb_pc=WB_reg_pc;


//***************    general register   ********************
wire [63:0] gpr[31:0];
wire [4:0]gpr_rd;
wire [63:0]gpr_wdata;
wire gpr_wen;

assign gpr_wen =  (reg_wr_ID == 5'b0)? 1'b0 : reg_wr_wen ;
assign gpr_rd  =  reg_wr_ID  ;
assign gpr_wdata = reg_wr_value ;

ysyx_22050612_RegisterFile #(5,64) cpu_gpr_group (clk, gpr_wdata, gpr_rd, gpr_wen, gpr);
//assign wen_fix = ( (rd != 5'b0)&&(exu_block == 1'b0) )?  wen : 1'b0;

reg [31:0]gpr_busy;
wire wen;
always@(posedge clk) begin
	if(rst) begin
		gpr_busy <= 32'b0;
	end
	if(gpr_rd != 5'b0 && gpr_wen == 1'b1 ) begin
		gpr_busy[gpr_rd] <= 1'b0;
	end
	if(rd != 5'b0 && wen == 1'b1 && ready_IF_ID == 1'b1 ) begin
		gpr_busy[rd]     <= 1'b1;
	end
end




//***************    control status register   ********************

wire [63:0]wdata_mtvec,wdata_mepc,wdata_mcause,wdata_mstatus;
wire [63:0]mtvec,mepc,mcause,mstatus;
wire wen_mtvec,wen_mepc,wen_mcause,wen_mstatus;
wire [63:0]src_csr;

//control and status register
ysyx_22050612_Reg #(64,64'h0) mtvec_csr           (clk, rst, wdata_mtvec  , mtvec  , wen_mtvec  );
ysyx_22050612_Reg #(64,64'h0) mepc_csr            (clk, rst, wdata_mepc   , mepc   , wen_mepc   );
ysyx_22050612_Reg #(64,64'h0) mcause_csr          (clk, rst, wdata_mcause , mcause , wen_mcause );
ysyx_22050612_Reg #(64,64'ha00001800) mstatus_csr (clk, rst, wdata_mstatus, mstatus, wen_mstatus);


//**************        processor       *******************
ysyx_22050612_IFU ifu (clk, rst, dnpc,valid_IF_ID, ready_IF_ID, pc_IF_ID, pc_update, inst_IF_ID , branch_flush);

wire       valid_IF_ID;
wire       ready_IF_ID;
wire [63:0]pc_IF_ID  ;
wire [31:0]inst_IF_ID;
assign pc = pc_IF_ID;

wire branch_flush;

ysyx_22050612_IDU idu (clk, rst, gpr, valid_IF_ID, ready_IF_ID, pc_IF_ID, inst_IF_ID, gpr_busy, mtvec, mepc, mcause, mstatus, /*imm_I,imm_U,imm_J,imm_B,imm_S,shamt, rd, rs1, rs2,*/ src_A,src_B, imm, rd, wen, opcode_ID_EX, valid_ID_EX, ready_ID_EX, pc_ID_EX, inst_ID_EX , EX_reg_valid,EX_reg_inst  , branch_flush);

wire       valid_ID_EX  ;
wire       ready_ID_EX  ;
wire [63:0]pc_ID_EX  ;
wire [31:0]inst_ID_EX;
wire [63:0]src_A;
wire [63:0]src_B;
wire [63:0]imm;
wire [23:0]opcode_ID_EX;
//wire [ 7:0]ALU_mode      ;
//wire [ 4:0]rd            ;


wire       EX_reg_valid;
wire [31:0]EX_reg_inst ;


ysyx_22050612_EXU exu (clk,rst, valid_ID_EX, ready_ID_EX, pc_ID_EX, inst_ID_EX,/*imm_I,imm_U,imm_J,imm_B,imm_S,shamt,rd,rs1,rs2,*/opcode_ID_EX,src_A,src_B,/*ALU_mode, src2, rd,*/ imm, dnpc,pc_update, valid_EX_MEM, ready_EX_MEM, pc_EX_MEM, inst_EX_MEM, opcode_EX_MEM, ALUoutput_EX_MEM , src_B_EX_MEM,/*reg_wr_wen, reg_wr_ID, reg_wr_value, */wdata_mtvec,wdata_mepc,wdata_mcause,wdata_mstatus,wen_mtvec,wen_mepc,wen_mcause,wen_mstatus,gpr , EX_reg_valid,EX_reg_inst,  MEM_reg_valid, MEM_reg_inst, MEM_reg_aluoutput, WB_reg_valid, WB_reg_inst, WB_reg_wdata  , branch_flush );

wire       valid_EX_MEM  ;
wire       ready_EX_MEM  ;
wire [63:0]pc_EX_MEM  ;
wire [31:0]inst_EX_MEM;
wire [23:0]opcode_EX_MEM;
wire [63:0]src_B_EX_MEM  ;
wire [63:0]ALUoutput_EX_MEM  ;

wire       MEM_reg_valid;
wire [31:0]MEM_reg_inst ;
wire [63:0]MEM_reg_aluoutput ;

ysyx_22050612_MEM mem (clk,rst, valid_EX_MEM, ready_EX_MEM, pc_EX_MEM, inst_EX_MEM,opcode_EX_MEM, ALUoutput_EX_MEM, src_B_EX_MEM, valid_MEM_WB, ready_MEM_WB, pc_MEM_WB, inst_MEM_WB, reg_wr_wen, reg_wr_ID, reg_wr_value,  MEM_reg_valid, MEM_reg_inst, MEM_reg_aluoutput , WB_reg_valid, WB_reg_inst, WB_reg_wdata);


wire       valid_MEM_WB  ;
wire       ready_MEM_WB  ;
wire [63:0]pc_MEM_WB  ;
wire [31:0]inst_MEM_WB;
wire       reg_wr_wen   ;
wire [ 4:0]reg_wr_ID    ;
wire [63:0]reg_wr_value ;

wire       WB_reg_valid;
wire [31:0]WB_reg_inst ;
wire [63:0]WB_reg_wdata ;

wire [63:0]WB_reg_pc ;

ysyx_22050612_WBU wbu (clk,rst, valid_MEM_WB, ready_MEM_WB, pc_MEM_WB, inst_MEM_WB, reg_wr_wen, reg_wr_ID, reg_wr_value, gpr , WB_reg_valid, WB_reg_inst, WB_reg_wdata, WB_reg_pc);





//************************  pipeline  ******************************

always @(negedge clk) begin
	//$display("busy %x",gpr_busy);
end

//*****************************************************************






/*
//*******************  axi  *******************************
wire arvalid_pc      ;  
wire [31:0]araddr_pc ;  
wire arready_pc      ;  
wire rvalid_pc       ;   
wire [63:0]rdata_pc  ; 
wire [1:0]rresp_pc   ;
wire rready_pc       ;

wire awvalid_pc      ;  
wire [31:0]awaddr_pc ; 
wire awready_pc      ; 
wire wvalid_pc       ;    
wire [63:0]wdata_pc  ;  
wire [7:0]wstrb_pc  ;  
wire wready_pc       ;      
wire [1:0]bresp_pc   ; 
wire bvalid_pc       ;   
wire bready_pc       ;   


wire arvalid_lsu      ;  
wire [31:0]araddr_lsu ;  
wire arready_lsu      ;  
wire rvalid_lsu       ;   
wire [63:0]rdata_lsu  ; 
wire [1:0]rresp_lsu   ;
wire rready_lsu       ;
wire awvalid_lsu      ;  
wire [31:0]awaddr_lsu ; 
wire awready_lsu      ; 
wire wvalid_lsu       ;    
wire [63:0]wdata_lsu  ;  
wire [7:0]wstrb_lsu  ;  
wire wready_lsu       ;      
wire [1:0]bresp_lsu   ; 
wire bvalid_lsu       ;   
wire bready_lsu       ;   


wire arvalid      ;  
wire [31:0]araddr ;  
wire arready      ;  
wire rvalid       ;   
wire [63:0]rdata  ; 
wire [1:0]rresp   ;
wire rready       ;
wire awvalid      ;  
wire [31:0]awaddr ; 
wire awready      ; 
wire wvalid       ;    
wire [63:0]wdata  ;  
wire [7:0]wstrb   ;  
wire wready       ;      
wire [1:0]bresp   ; 
wire bvalid       ;   
wire bready       ;  



//ysyx_22050612_SRAM sram_pc (clk,rst,arvalid_pc,araddr_pc,arready_pc,rvalid_pc,rdata_pc,rresp_pc,rready_pc, 1'b0, 32'b0,  , 1'b0, 64'b0, 8'b0, , , , 1'b0);
//ysyx_22050612_SRAM sram_pc (clk,rst,arvalid_pc,araddr_pc,arready_pc,rvalid_pc,rdata_pc,rresp_pc,rready_pc,awvalid_pc,awaddr_pc,awready_pc,wvalid_pc,wdata_pc,wstrb_pc,wready_pc,bresp_pc,bvalid_pc,bready_pc);

//ysyx_22050612_SRAM sram (clk,rst,arvalid_lsu,araddr_lsu,arready_lsu,rvalid_lsu,rdata_lsu,rresp_lsu,rready_lsu,awvalid_lsu,awaddr_lsu,awready_lsu,wvalid_lsu,wdata_lsu,wstrb_lsu,wready_lsu,bresp_lsu,bvalid_lsu,bready_lsu);
ysyx_22050612_SRAM sram (clk,rst,arvalid,araddr,arready,rvalid,rdata,rresp,rready,awvalid,awaddr,awready,wvalid,wdata,wstrb,wready,bresp,bvalid,bready);

ysyx_22050612_Arbiter arbiter (clk,rst,
	arvalid_pc,arvalid_lsu,arvalid,
	araddr_pc,araddr_lsu,araddr,
	arready_pc,arready_lsu,arready,
	rvalid_pc,rvalid_lsu,rvalid,
	rdata_pc,rdata_lsu,rdata,
	rresp_pc,rresp_lsu,rresp,
	rready_pc,rready_lsu,rready,
	awvalid_pc,awvalid_lsu,awvalid,
	awaddr_pc,awaddr_lsu,awaddr,
	awready_pc,awready_lsu,awready,
	wvalid_pc,wvalid_lsu,wvalid,
	wdata_pc,wdata_lsu,wdata,
	wstrb_pc,wstrb_lsu,wstrb,
	wready_pc,wready_lsu,wready,
	bresp_pc,bresp_lsu,bresp,
	bvalid_pc,bvalid_lsu,bvalid,
	bready_pc,bready_lsu,bready);
//	1'b0,awvalid_lsu,awvalid,
//	32'b0,awaddr_lsu,awaddr,
//	1'b0,awready_lsu,awready,
//	1'b0,wvalid_lsu,wvalid,
//	64'b0,wdata_lsu,wdata,
//	8'b0,wstrb_lsu,wstrb,
//	1'b0,wready_lsu,wready,
//	2'b0,bresp_lsu,bresp,
//	1'b0,bvalid_lsu,bvalid,
//	1'b0,bready_lsu,bready);

//************************************************************
*/



//always @(posedge clk) begin
//  $display("%x",inst);
//end

initial set_gpr_ptr(gpr); 

endmodule
