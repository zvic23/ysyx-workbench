module ysyx_22050612_IDU(
input [31:0]inst;




output imm,
output opcode


);







endmodule
