module ysyx_22050612_IDU(
input clk,
input [31:0]inst,




output [63:0]imm_I,
output [ 4:0]rd,
output [ 4:0]rs1,
output [ 4:0]rs2,
output [ 2:0]opcode


);

assign rd = inst[11: 7];
assign rs1= inst[19:15];
assign rs2= inst[24:20];

assign imm_I= (inst[31]==1'b1)?{{52{1'b1}},inst[31:20]}:{{52{1'b0}},inst[31:20]};

ysyx_22050612_MuxKey #(1, 3, 3) a3 (opcode, inst[2:0], {
    3'b011, 3'b1
  });

  always @(posedge clk) begin
    $display("%x,%d",inst,opcode);
  end





endmodule
